module test_tb();
reg clk;
reg[8192:0] s;
//----------------
wire[9209:0] c;
//-----------------
test u1(
.clk(clk),
.s(s),
.c(c)
);
//------------------------------------------
task Loading;
begin
	  s[8192:7590] <= 603'O2_3_3_4_6_1_6_6_2_3_4_5_5_5_3_3_7_4_6_2_4_4_7_1_4_4_1_6_6_3_5_1_4_2_3_6_1_2_3_2_6_7_1_2_5_3_7_7_5_6_3_4_7_4_7_5_3_4_6_1_3_7_3_5_6_7_5_1_0_4_4_7_5_5_4_2_7_4_0_5_4_0_6_2_2_1_2_2_5_0_2_2_6_3_5_4_5_1_7_6_0_3_2_4_2_4_4_4_3_0_4_3_1_3_3_4_6_5_6_0_2_3_7_6_3_2_0_5_4_1_3_1_5_3_7_0_6_4_4_5_5_1_6_0_2_1_6_0_4_4_5_6_0_6_4_5_1_4_5_7_3_1_0_4_6_5_2_7_4_7_1_1_5_6_5_2_1_6_5_2_2_2_6_6_4_4_2_5_6_3_3_3_2_5_6_6_5_2_5_1_1;
    s[7589:6990] <= 600'O1_1_4_1_6_5_6_3_5_6_4_2_7_0_2_7_3_2_1_6_1_2_6_3_4_4_5_0_4_0_6_2_6_2_4_7_0_0_0_5_4_1_6_4_0_0_1_6_1_2_2_1_6_5_5_5_4_2_5_1_1_0_7_7_1_3_5_2_5_4_3_2_5_6_5_3_7_2_4_7_2_2_6_0_2_4_1_4_6_4_5_6_2_4_1_4_6_6_3_2_5_6_4_7_1_1_2_3_3_2_5_1_3_2_2_1_4_2_1_0_2_4_6_0_6_1_6_6_6_1_4_3_1_4_4_2_4_7_3_5_3_0_2_6_2_1_4_3_5_4_6_6_1_1_6_4_0_6_4_4_4_5_6_3_1_5_2_6_3_6_1_1_6_0_5_5_3_3_7_3_3_1_2_2_6_2_2_3_5_1_6_1_3_0_5_5_2_5_4_6;
    s[6989:6390] <= 600'O4_6_3_3_3_2_7_3_2_3_5_3_1_6_4_3_2_2_4_3_5_0_6_5_1_6_1_4_4_1_0_5_5_3_0_4_1_5_4_2_6_5_6_0_1_5_5_5_4_3_4_6_5_4_2_5_3_4_6_6_6_7_6_0_0_1_2_0_3_2_4_6_2_2_6_2_1_4_6_3_5_4_3_3_7_1_2_3_4_6_3_3_5_3_6_3_3_3_2_1_0_6_2_6_5_6_7_1_3_7_5_6_3_0_4_2_4_5_4_4_3_2_3_0_4_7_1_0_6_2_0_6_1_6_1_2_4_4_5_5_3_1_5_2_5_6_1_7_0_6_6_0_4_7_2_6_4_6_6_0_2_5_3_7_5_4_2_2_6_3_6_1_6_0_6_6_4_1_1_5_6_0_5_7_2_4_2_2_6_5_2_4_3_1_0_3_2_2_2_1;
    s[6389:5790] <= 600'O3_5_1_5_3_3_1_1_4_2_4_7_5_5_7_5_4_7_0_2_7_5_3_5_3_3_1_3_0_3_2_7_4_6_3_3_6_7_4_6_5_4_7_6_7_5_3_3_6_0_1_3_4_0_5_6_1_3_2_7_4_2_1_4_6_6_6_1_4_6_1_6_6_2_1_3_6_3_3_4_1_1_6_4_2_6_0_3_5_2_3_4_6_5_0_2_3_6_3_2_4_3_6_7_6_5_5_6_0_2_0_6_4_3_2_4_2_0_1_0_3_1_3_6_2_1_4_6_2_0_1_1_5_3_5_5_4_4_6_5_6_3_1_0_5_2_5_5_4_5_4_3_3_7_3_1_2_5_6_7_2_5_4_3_4_3_5_5_2_1_6_3_5_1_1_6_6_7_6_0_4_7_4_6_0_7_6_4_3_2_5_0_3_6_4_3_3_2_7_7;
    s[5789:5190] <= 600'O4_7_3_3_1_1_6_5_4_6_4_4_1_4_1_0_5_4_2_3_4_4_1_1_0_3_3_1_5_0_1_7_7_0_3_6_2_6_6_4_0_3_6_5_3_4_2_4_7_6_2_5_3_7_1_2_6_1_4_6_5_1_3_2_3_4_1_6_4_1_4_7_5_5_3_2_4_2_2_6_6_6_6_1_4_4_6_5_3_5_6_4_1_6_0_4_1_3_6_2_6_5_3_2_2_5_0_5_4_5_7_3_2_6_6_3_1_4_1_4_2_2_5_4_6_1_5_0_6_5_7_1_6_4_4_2_1_6_1_3_4_7_4_7_2_3_5_0_5_3_6_3_2_7_5_3_1_5_4_1_1_7_3_0_0_1_6_3_4_3_0_6_2_2_4_3_3_5_7_4_2_1_3_0_6_4_1_4_0_6_3_4_4_5_3_1_3_0_5_0;
    s[5189:4590] <= 600'O7_5_7_4_2_2_5_7_2_5_1_4_3_5_2_1_3_4_1_3_5_6_2_3_6_5_2_5_2_2_0_3_3_2_2_2_7_6_3_3_4_3_2_7_1_6_0_2_5_5_1_7_4_2_4_6_6_3_3_2_0_5_1_2_3_6_0_6_2_2_3_5_1_2_7_4_2_7_6_1_0_5_6_1_0_4_4_4_0_5_7_6_1_2_2_4_4_2_6_6_5_2_0_5_7_1_1_6_3_6_6_1_2_0_4_5_4_0_7_4_2_1_4_4_5_1_2_1_6_2_2_0_6_3_4_6_5_5_1_4_7_4_6_7_6_1_0_3_0_3_7_2_3_3_6_6_3_3_6_5_5_7_4_6_3_6_3_5_7_4_3_1_2_1_3_2_2_6_4_4_5_1_4_2_2_4_6_1_5_6_1_2_3_6_4_2_4_4_3_0;
    s[4589:3990] <= 600'O5_4_3_0_3_2_1_6_3_0_3_5_1_6_2_2_1_5_0_7_1_2_5_1_4_5_7_5_5_3_2_4_2_6_5_6_6_3_2_5_7_5_6_5_4_5_3_6_0_7_1_4_3_1_5_4_5_4_6_4_7_6_4_6_3_6_2_7_2_1_5_6_6_2_6_4_3_6_7_1_5_2_3_2_6_7_5_5_7_5_4_3_4_3_3_3_3_4_6_1_2_4_3_2_4_6_0_3_1_4_4_5_2_4_3_6_5_2_2_2_7_2_1_3_5_5_5_0_3_6_2_4_2_1_3_6_7_6_1_2_2_2_7_4_5_6_1_6_1_5_5_5_1_3_4_4_6_5_6_4_7_0_4_2_3_5_1_4_2_6_1_1_7_1_1_1_1_3_5_6_6_5_3_5_7_4_2_6_2_2_3_4_4_1_1_2_5_3_6_7;
    s[3989:3390] <= 600'O3_0_4_5_2_3_2_7_3_4_2_1_0_6_5_1_6_5_5_7_0_3_3_4_1_5_0_4_5_3_4_1_5_3_1_3_2_2_4_4_3_2_6_6_2_4_5_7_6_3_1_6_1_1_2_6_4_4_6_4_0_6_4_3_2_2_3_2_0_1_2_1_4_6_6_6_5_6_5_1_7_1_5_2_2_2_1_4_7_3_4_4_5_3_6_6_5_2_6_1_4_4_5_3_5_6_0_1_6_3_3_7_5_7_2_1_3_4_4_7_3_3_7_2_5_7_5_2_4_0_6_3_2_7_3_2_1_4_1_1_4_2_3_5_6_2_7_7_1_5_4_6_4_5_5_3_2_0_3_5_2_4_2_2_5_6_6_1_3_6_2_7_4_1_6_5_4_2_0_2_3_4_7_1_5_6_3_1_6_3_1_6_4_1_6_0_0_7_5_3;
    s[3389:2790] <= 600'O4_5_0_5_5_3_4_2_1_3_6_2_3_2_1_4_6_6_5_3_2_5_6_6_1_3_1_2_6_1_1_4_2_3_6_6_5_3_5_1_4_5_4_2_3_1_6_3_2_5_2_6_6_6_3_3_6_3_4_5_7_4_4_4_6_6_1_1_2_5_1_7_5_1_6_6_7_4_4_1_4_4_1_3_4_1_4_0_2_4_2_4_3_1_6_4_5_5_5_6_4_1_3_6_1_2_7_6_2_7_0_3_3_3_1_3_4_7_2_2_2_2_1_0_3_2_6_4_6_7_4_1_6_4_6_3_4_0_6_4_1_5_3_1_2_2_2_5_5_4_4_4_7_4_4_6_4_2_7_3_4_5_5_1_1_2_6_4_3_3_5_5_5_1_3_4_3_3_2_5_3_5_3_5_7_4_6_2_6_1_3_0_6_1_1_1_5_1_2_5;
    s[2789:2190] <= 600'O4_6_0_3_4_4_6_1_2_0_7_5_5_1_2_1_3_6_4_5_4_5_6_4_1_4_1_6_1_2_4_3_6_4_2_5_1_5_4_2_1_1_1_1_7_0_7_0_7_2_4_6_6_1_5_7_7_1_1_5_0_0_3_6_7_0_4_6_6_6_6_5_1_4_1_6_6_1_6_3_3_2_6_5_3_5_7_1_2_4_6_6_3_1_1_3_6_2_6_5_0_6_6_3_6_1_5_6_6_2_1_4_3_3_7_4_7_3_3_5_5_3_0_1_6_5_0_4_5_1_2_6_1_6_6_0_3_1_4_1_0_7_7_3_5_0_1_0_3_1_7_3_7_5_4_4_5_0_5_6_0_6_5_7_2_6_4_1_2_5_6_1_3_2_6_2_6_2_6_1_5_0_4_4_3_1_6_1_3_0_1_3_6_1_5_5_0_3_7_1;
    s[2189:1590] <= 600'O5_4_4_3_4_3_1_2_4_4_7_7_1_5_4_3_2_3_5_7_1_6_4_6_1_2_0_4_5_2_2_2_3_5_4_3_6_7_4_1_4_3_7_2_5_4_1_5_0_1_0_6_6_1_3_1_4_7_2_7_2_1_5_7_4_0_3_1_2_0_6_6_3_6_5_4_3_3_1_2_4_3_5_4_6_1_3_4_1_4_0_4_6_3_3_1_0_5_6_2_1_3_6_6_5_7_7_1_5_3_0_6_3_5_0_2_5_1_4_3_5_5_3_2_2_6_3_3_3_7_2_6_0_2_5_2_4_3_0_4_4_5_2_3_5_6_0_1_5_5_7_1_3_5_3_6_2_1_5_1_6_5_3_0_1_2_6_4_2_2_3_6_6_4_4_5_0_4_0_3_3_0_0_6_4_3_3_1_1_2_2_5_3_3_1_6_5_6_5_7;
    s[1589: 990] <= 600'O7_2_4_5_3_6_1_1_0_1_4_4_3_2_0_6_4_3_2_6_6_6_3_7_6_1_2_6_3_3_7_7_5_4_6_3_1_2_2_4_0_0_1_7_6_5_7_7_7_1_7_4_1_2_6_6_0_4_6_2_0_2_1_3_3_3_6_3_2_0_2_2_0_5_0_4_3_2_5_2_1_4_1_6_5_6_5_6_4_5_5_2_4_6_0_4_3_6_4_7_4_6_3_4_1_4_7_4_3_6_1_6_0_4_5_4_3_2_4_6_5_7_1_4_1_4_5_1_5_3_6_2_0_2_1_7_0_1_0_2_0_4_4_2_1_1_3_0_4_3_2_5_6_2_4_3_2_6_7_4_1_1_4_2_2_4_1_5_0_0_2_1_6_6_3_1_3_3_5_3_7_6_7_2_2_6_1_1_4_6_3_2_1_7_4_3_5_6_2_5;
    s[ 989: 390] <= 600'O1_7_5_1_3_4_7_4_4_5_6_1_3_2_5_6_3_6_2_4_3_6_5_6_1_2_5_2_0_3_7_2_4_3_0_4_6_2_0_2_5_2_5_0_5_3_0_3_5_6_7_7_6_6_6_4_3_1_5_6_2_6_0_3_2_1_4_2_7_3_5_0_4_4_6_5_6_6_1_1_6_0_3_2_5_1_6_5_4_2_0_4_0_0_1_3_5_6_3_0_2_4_6_2_3_6_4_4_2_3_6_2_3_3_5_4_5_3_3_3_0_3_7_5_5_5_5_6_5_7_1_3_3_2_0_7_5_1_1_5_3_1_3_1_6_7_0_5_5_2_6_2_0_1_6_5_5_4_6_0_3_2_3_6_2_4_0_1_6_1_6_2_5_0_5_3_7_2_3_1_7_3_1_5_4_2_5_6_2_4_3_1_4_7_1_6_4_3_1_2;
    s[ 389:   0] <= 600'O3_4_2_5_6_5_3_4_4_1_3_2_4_7_3_0_7_6_3_2_6_4_4_5_1_6_7_1_6_6_0_4_5_3_5_5_4_4_2_6_3_4_6_2_3_4_3_1_5_0_3_0_7_4_6_3_6_2_6_6_3_4_4_6_1_0_6_2_2_4_2_6_6_7_3_6_1_4_5_1_4_6_2_2_6_3_1_2_5_4_2_4_5_2_3_3_5_1_6_2_3_5_5_1_5_1_7_6_4_5_7_1_5_6_5_1_3_0_2_1_3_4_6_3_4_6_6_4_6_0;
    $display("Loading is successful!!!!");
end
endtask
//-------------------------------
initial begin
	  clk = 1'b0;
	  Loading;
#10
    clk = 1'b1;
#10
    clk = 1'b0;

    $display("the c is %O %O %O %O %O %O %O %O %O %O %O %O %O %O %O %O %O %O %O %O",
    c[59:57],c[56:54],c[53:51],c[50:48],c[47:45],c[44:42],c[41:39],c[38:36],c[35:33],c[32:30],
    c[29:27],c[26:24],c[23:21],c[20:18],c[17:15],c[14:12],c[11:9],c[8:6],c[5:3],c[2:0]);
end
endmodule

